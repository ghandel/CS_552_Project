module and4 (A, B, C, D, out);

    input A;
    input B;
    input C;
    input D;
    
    output out;
    
    assign out = A & B & C & D;

endmodule
